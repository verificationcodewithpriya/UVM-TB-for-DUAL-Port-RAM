package env_pkg;
 import uvm_pkg :: *;
`include "uvm_macros.svh"

`include "config_obj.sv"
`include "transaction.sv"
`include "seq.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "func_cvg.sv"
`include "environment.sv"
`include "test.sv"

endpackage

